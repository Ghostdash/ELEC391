module LFSR (
  input logic clk,
  output logic [7:0] lfsr_out
);

  logic [7:0] lfsr_reg=8'b10000001;  
  logic feedback;

  always @(posedge clk) begin
     lfsr_reg <= {lfsr_reg[6:0], feedback};
  end

  assign feedback = lfsr_reg[7] ^ lfsr_reg[5] ^ lfsr_reg[4] ^ lfsr_reg[3];

  assign lfsr_out = lfsr_reg;

endmodule 