module QAM16 ();
    



endmodule