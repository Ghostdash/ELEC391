module tb_qpsk_hamming();
    logic clk, reset;
    

    Hamming_encoder encoder();
    Hamming_decoder decoder();
    QPSK_mod modulator();
    QPSK_demod demodulator();





endmodule